module hello_module;

initial begin
        $display("Hello, world!");
        $finish();
        end

endmodule
