module hello_module;

initial begin
        $display("Hello, world!", magic);
        $finish();
        end

endmodule
