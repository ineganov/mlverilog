module Blah(a,b,c);
  
    input [1:0] a,wert, khkhhkhkhkhk_h;
    input b;
    wire dsfgsdfg;
    reg h,j,k;

    pqpq instance_name1 (.x(a),
                         .y(b) ) ;

    pqpq # (.QWE(RTY)) instance_name2 ( .x(a),
                         .y({a,b,3+2}) ) ;

    assign a = b;
    assign {q,w,e} = 4+1;

endmodule